version https://git-lfs.github.com/spec/v1
oid sha256:8731c07e320af08e3f24afec59739dab22f87bc6363bfdc5fdbefb9e941d9785
size 104858112
